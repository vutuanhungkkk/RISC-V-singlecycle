module decoder(
   input clk,
	input [31:0] instr,
	output [4:0] rd_addr,
	output [4:0] rs1_addr,
	output [4:0] rs2_addr
	);

	assign rs1_addr = instr[19:15];
	assign rs2_addr = instr[24:20];
	assign rd_addr = instr[11:7];

endmodule