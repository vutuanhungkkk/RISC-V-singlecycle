// Module to generate immediate values based on instruction type
module ImmGen(
    input wire [31:0] instr, // 32-bit instruction input
    output reg [31:0] Imm // 32-bit immediate output
);

    wire [4:0] srai;
    assign srai = instr[24:20]; // Extract bits 24:20 for SRAI immediate
    always @(*) begin
        case(instr[6:0])
            // I-type load instructions
            7'b0000011: Imm = {instr[31] ? {20{1'b1}} : 20'b0, instr[31:20]};
            // I-type addi instructions
            7'b0010011: begin
                // Check for SRAI, SLLI, and SRLI instructions
                if ((instr[31:25] == 7'b0100000 && instr[14:12] == 3'b101) ||
                    (instr[14:12] == 3'b001) || (instr[14:12] == 3'b101)) begin
                    // Set immediate value based on srai
                    Imm = {srai[4] ? {27{1'b1}} : 27'b0, srai};
                end else begin
                    // Otherwise, set immediate value based on bits 31:20
                    Imm = {instr[31] ? {20{1'b1}} : 20'b0, instr[31:20]};
                end
            end

            // S-type store instructions
            7'b0100011: Imm = {instr[31] ? {20{1'b1}} : 20'b0, instr[31:25], instr[11:7]};

            // B-type branch instructions
            7'b1100011: Imm = {instr[31] ? {20{1'b1}} : 20'b0, instr[7], instr[30:25], instr[11:8], 1'b0};

            // JALR instructions
            7'b1100111: Imm = {instr[31] ? {20{1'b1}} : 20'b0, instr[30:25], instr[24:21], instr[20]};

            // U-type instructions (LUI and AUIPC)
            7'b0010111, 7'b0110111: Imm = {instr[31:12], 12'b0};

            // JAL instructions
            7'b1101111: Imm = {instr[31] ? {20{1'b1}} : 20'b0, instr[19:12], instr[19:12], instr[20], instr[30:25], instr[24:21], 1'b0};
            default: 
                Imm = 32'b0;
        endcase
    end
endmodule
